library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity LOAD_BALANCER is
	PORT (
			CORE_ID 	: IN STD_LOGIC;
			
			ADDRESS_A_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_B_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_C_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_0_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_1_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_W_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			DATA_TO_W_C0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			W_EN_C0		  : IN STD_LOGIC;
			
			ADDRESS_A_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_B_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_C_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_0_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_1_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_W_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			DATA_TO_W_C1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			W_EN_C1		  : IN STD_LOGIC;
			
			ADDRESS_IO		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			DATA_IO			: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			IO_ENABLE		: IN STD_LOGIC;
			
			global_enable	: IN STD_LOGIC_VECTOR (5 downto 0);

			ADDRESS_A_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_B_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_C_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_0_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_1_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			ADDRESS_W_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			DATA_TO_W_MAG  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			W_EN_MAG		  	: OUT STD_LOGIC

			);
end;

architecture balancer of LOAD_BALANCER is
	
begin
	
	process (CORE_ID, ADDRESS_A_C0, ADDRESS_B_C0, ADDRESS_C_C0, ADDRESS_0_C0, ADDRESS_1_C0, ADDRESS_W_C0, 
				ADDRESS_A_C1, ADDRESS_B_C1, ADDRESS_C_C1, ADDRESS_0_C1, ADDRESS_1_C1, ADDRESS_W_C1,
				DATA_TO_W_C0, DATA_TO_W_C1, W_EN_C0, W_EN_C1, IO_ENABLE, ADDRESS_IO, DATA_IO, global_enable) begin
		if (CORE_ID = '0') then
			if (IO_ENABLE = '1') then
				ADDRESS_A_MAG <= "00000000000000000000000000000000";
				ADDRESS_B_MAG <= "00000000000000000000000000000001";
				ADDRESS_C_MAG <= "00000000000000000000000000000010";
				ADDRESS_0_MAG <= "00000000000000000000000000000011";
				ADDRESS_1_MAG <= "00000000000000000000000000000100";
				DATA_TO_W_MAG <= DATA_IO;
				ADDRESS_W_MAG <= ADDRESS_IO;
				W_EN_MAG <= '1';
			else
				ADDRESS_A_MAG <= ADDRESS_A_C0;
				ADDRESS_B_MAG <= ADDRESS_B_C0;
				ADDRESS_C_MAG <= ADDRESS_C_C0;
				ADDRESS_0_MAG <= ADDRESS_0_C0;
				ADDRESS_1_MAG <= ADDRESS_1_C0;
				ADDRESS_W_MAG <= ADDRESS_W_C0;
				DATA_TO_W_MAG <= DATA_TO_W_C0;
				W_EN_MAG <= W_EN_C0;
			end if;
		else
			if (IO_ENABLE = '1') then
				ADDRESS_A_MAG <= "00000000000000000000000000000000";
				ADDRESS_B_MAG <= "00000000000000000000000000000001";
				ADDRESS_C_MAG <= "00000000000000000000000000000010";
				ADDRESS_0_MAG <= "00000000000000000000000000000011";
				ADDRESS_1_MAG <= "00000000000000000000000000000100";
				DATA_TO_W_MAG <= DATA_IO;
				ADDRESS_W_MAG <= ADDRESS_IO;
				W_EN_MAG <= '1';
			else
				ADDRESS_A_MAG <= ADDRESS_A_C1;
				ADDRESS_B_MAG <= ADDRESS_B_C1;
				ADDRESS_C_MAG <= ADDRESS_C_C1;
				ADDRESS_0_MAG <= ADDRESS_0_C1;
				ADDRESS_1_MAG <= ADDRESS_1_C1;
				ADDRESS_W_MAG <= ADDRESS_W_C1;
				DATA_TO_W_MAG <= DATA_TO_W_C1;
				W_EN_MAG <= W_EN_C1;
			end if;
		end if;
	end process;

end;