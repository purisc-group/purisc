library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MAGIC_tb is
end;

architecture testing of MAGIC_tb is
	component MAGIC
		PORT (
				ADDRESS_A  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				ADDRESS_B  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				ADDRESS_C  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				ADDRESS_0  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				ADDRESS_1  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				ADDRESS_W  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				DATA_TO_W  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
				W_EN		  : IN STD_LOGIC;
				CLK		  : IN STD_LOGIC;
				RESET_n    : IN STD_LOGIC;
				DATA_OUT_A : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				DATA_OUT_B : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				DATA_OUT_C : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				DATA_OUT_0 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				DATA_OUT_1 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				STALL		  : OUT STD_LOGIC
				);
	end component;
	
	signal ADDRESS_A  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal ADDRESS_B  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal ADDRESS_C  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal ADDRESS_0  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal ADDRESS_1  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal ADDRESS_W  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal DATA_TO_W  : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal W_EN		  : STD_LOGIC := '0';
	signal CLK		  : STD_LOGIC := '1';
	signal RESET_n    : STD_LOGIC := '0';
	signal DATA_OUT_A : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal DATA_OUT_B : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal DATA_OUT_C : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal DATA_OUT_0 : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal DATA_OUT_1 : STD_LOGIC_VECTOR (31 DOWNTO 0);
	signal STALL		  : STD_LOGIC;
	
	constant clk_period : time := 10ns;
	
begin

	uut : MAGIC PORT MAP (
								ADDRESS_A,
								ADDRESS_B,
								ADDRESS_C,
								ADDRESS_0,
								ADDRESS_1,
								ADDRESS_W,
								DATA_TO_W,
								W_EN,
								CLK,
								RESET_n,
								DATA_OUT_A,
								DATA_OUT_B,
								DATA_OUT_C,
								DATA_OUT_0,
								DATA_OUT_1,
								STALL
								);
	
	clk_process : process begin
		clk <= '1';
		wait for clk_period/2;
		clk <= '0';
		wait for clk_period/2;
	end process;
	
	stim_process : process begin
		wait for 20 ns;
		ADDRESS_A <= "00000000000000000000000000000000";
		ADDRESS_B <= "00000000000000000000000000000001";
		ADDRESS_C <= "00000000000000000000000000000010";
		ADDRESS_0 <= "00000000000000000000000000000011";
		ADDRESS_1 <= "00000000000000000000000000000100";
		RESET_n <= '1';
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000000";
		DATA_TO_W <= "00000000000000000000000000000000";
		W_EN <= '1';
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000001";
		DATA_TO_W <= "00000000000000000000000000000001";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000010";
		DATA_TO_W <= "00000000000000000000000000000010";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000011";
		DATA_TO_W <= "00000000000000000000000000000011";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000100";
		DATA_TO_W <= "00000000000000000000000000000100";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000101";
		DATA_TO_W <= "00000000000000000000000000000101";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000110";
		DATA_TO_W <= "00000000000000000000000000000110";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000000111";
		DATA_TO_W <= "00000000000000000000000000000111";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001000";
		DATA_TO_W <= "00000000000000000000000000001000";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001001";
		DATA_TO_W <= "00000000000000000000000000001001";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001010";
		DATA_TO_W <= "00000000000000000000000000001010";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001011";
		DATA_TO_W <= "00000000000000000000000000001011";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001100";
		DATA_TO_W <= "00000000000000000000000000001100";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001101";
		DATA_TO_W <= "00000000000000000000000000001101";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001110";
		DATA_TO_W <= "00000000000000000000000000001110";
		wait for clk_period;
		ADDRESS_W <= "00000000000000000000000000001111";
		DATA_TO_W <= "00000000000000000000000000001111";
		wait for clk_period;
		ADDRESS_A <= "00000000000000000000000000000110";
		ADDRESS_B <= "00000000000000000000000000001100";
		ADDRESS_C <= "00000000000000000000000000000111";
		ADDRESS_0 <= "00000000000000000000000000001000";
		ADDRESS_1 <= "00000000000000000000000000001001";
		W_EN <= '0';
		wait;
	end process;
end;